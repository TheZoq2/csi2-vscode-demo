module launder_clock(input clk_i, output clk_o, output output__);
    assign clk_o = clk_i;
endmodule
